library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sp0256_256b_019_decoded is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sp0256_256b_019_decoded is
	type rom is array(0 to  11295) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"18",X"01",X"00",X"19",X"01",X"00",X"1A",X"01",X"00",X"1B",X"01",X"00",X"1C",X"01",X"00",
		X"1D",X"0A",X"00",X"27",X"0A",X"00",X"31",X"01",X"00",X"32",X"03",X"00",X"35",X"03",X"00",X"38",
		X"03",X"00",X"3B",X"03",X"00",X"3E",X"01",X"00",X"3F",X"04",X"00",X"43",X"06",X"00",X"49",X"01",
		X"00",X"4A",X"04",X"00",X"4E",X"03",X"00",X"51",X"02",X"00",X"53",X"06",X"00",X"59",X"08",X"00",
		X"61",X"02",X"00",X"63",X"03",X"00",X"66",X"01",X"00",X"67",X"03",X"00",X"6A",X"06",X"00",X"70",
		X"01",X"00",X"71",X"03",X"00",X"74",X"02",X"00",X"76",X"01",X"00",X"77",X"01",X"00",X"78",X"03",
		X"00",X"7B",X"05",X"00",X"80",X"03",X"00",X"83",X"02",X"00",X"85",X"03",X"00",X"88",X"03",X"00",
		X"8B",X"03",X"00",X"8E",X"02",X"00",X"90",X"03",X"00",X"93",X"01",X"00",X"94",X"03",X"00",X"97",
		X"04",X"00",X"9B",X"03",X"00",X"9E",X"04",X"00",X"A2",X"03",X"00",X"A5",X"04",X"00",X"A9",X"0D",
		X"00",X"B6",X"04",X"00",X"BA",X"04",X"00",X"BE",X"03",X"00",X"C1",X"09",X"00",X"CA",X"0A",X"00",
		X"D4",X"07",X"00",X"DB",X"02",X"00",X"DD",X"01",X"00",X"DE",X"06",X"00",X"E4",X"03",X"00",X"E7",
		X"09",X"00",X"F0",X"09",X"00",X"F9",X"08",X"01",X"01",X"02",X"01",X"03",X"03",X"01",X"06",X"03",
		X"01",X"09",X"13",X"01",X"1C",X"16",X"01",X"32",X"12",X"01",X"44",X"1B",X"01",X"5F",X"19",X"01",
		X"78",X"1A",X"01",X"92",X"13",X"01",X"A5",X"0E",X"01",X"B3",X"16",X"01",X"C9",X"18",X"01",X"E1",
		X"1D",X"01",X"FE",X"01",X"01",X"FF",X"01",X"02",X"00",X"01",X"02",X"01",X"01",X"02",X"02",X"01",
		X"02",X"03",X"01",X"02",X"04",X"01",X"02",X"05",X"01",X"02",X"06",X"01",X"02",X"07",X"01",X"02",
		X"08",X"01",X"02",X"09",X"01",X"02",X"0A",X"01",X"02",X"0B",X"01",X"02",X"0C",X"01",X"02",X"0D",
		X"01",X"02",X"0E",X"01",X"02",X"0F",X"01",X"02",X"10",X"01",X"02",X"11",X"01",X"02",X"12",X"01",
		X"02",X"13",X"01",X"02",X"14",X"01",X"02",X"15",X"01",X"02",X"16",X"01",X"02",X"17",X"00",X"02",
		X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",
		X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",
		X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"00",X"02",X"17",X"0A",X"02",X"21",X"0C",X"02",
		X"2D",X"11",X"02",X"3E",X"10",X"02",X"4E",X"12",X"02",X"60",X"18",X"02",X"78",X"0F",X"02",X"87",
		X"1F",X"02",X"A6",X"18",X"02",X"BE",X"01",X"02",X"BF",X"01",X"02",X"C0",X"01",X"02",X"C1",X"01",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"01",X"40",X"5B",X"A0",X"60",X"B8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"00",X"C0",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"02",X"00",X"50",X"5B",X"A0",X"60",X"A8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"02",X"00",X"80",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"00",X"70",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"00",X"A0",X"5B",X"A0",X"60",X"B8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"04",X"01",X"C0",X"5B",X"A8",X"60",X"C0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"A8",X"60",X"D0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"04",X"02",X"80",X"5B",X"A8",X"60",X"E0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"09",X"01",X"00",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"03",X"00",X"5B",X"B0",X"70",X"C8",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"01",X"02",X"80",X"5B",X"C8",X"70",X"B0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"03",X"00",X"5B",X"C8",X"70",X"B0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"02",X"80",X"5B",X"B0",X"70",X"C8",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"02",X"00",X"5B",X"C8",X"70",X"F8",X"70",X"B8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"B0",X"70",X"D0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"03",X"03",X"80",X"5B",X"B0",X"70",X"F8",X"70",X"E0",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"03",X"00",X"5B",X"A8",X"70",X"E0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"A0",X"70",X"E8",X"70",X"00",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"03",X"01",X"00",X"5B",X"A0",X"70",X"F0",X"70",X"00",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"07",X"06",X"00",X"5B",X"00",X"50",X"28",X"50",X"40",X"50",X"F8",X"10",X"E8",X"58",X"AA",X"64",
		X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"40",X"FC",X"04",X"CB",X"68",
		X"07",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"20",X"40",X"C5",X"62",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"F4",X"2C",X"BF",X"3B",
		X"07",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"50",X"F8",X"44",X"CF",X"3A",
		X"05",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"18",X"42",X"FA",X"30",
		X"04",X"01",X"C0",X"5B",X"18",X"60",X"30",X"50",X"38",X"20",X"00",X"10",X"00",X"60",X"E6",X"38",
		X"05",X"01",X"40",X"5B",X"18",X"50",X"28",X"40",X"40",X"30",X"FC",X"68",X"E8",X"52",X"DD",X"16",
		X"04",X"00",X"E0",X"5B",X"00",X"30",X"18",X"20",X"38",X"40",X"FC",X"60",X"E0",X"2A",X"A1",X"54",
		X"03",X"01",X"40",X"5B",X"08",X"30",X"20",X"30",X"20",X"10",X"FC",X"68",X"E8",X"1C",X"A2",X"50",
		X"05",X"01",X"80",X"5B",X"08",X"30",X"20",X"40",X"20",X"10",X"FC",X"68",X"E0",X"24",X"9B",X"5B",
		X"06",X"06",X"00",X"5B",X"00",X"50",X"10",X"20",X"30",X"50",X"E8",X"60",X"34",X"1E",X"A0",X"6E",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"28",X"1C",X"4E",X"F4",X"21",
		X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"1C",X"44",X"EA",X"53",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"1C",X"46",X"E7",X"5A",
		X"06",X"00",X"1C",X"5B",X"98",X"60",X"C0",X"60",X"E0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"03",X"00",X"50",X"5B",X"98",X"60",X"C0",X"60",X"E8",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"01",X"00",X"C0",X"5B",X"98",X"60",X"C0",X"60",X"E8",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"02",X"02",X"80",X"5B",X"A0",X"60",X"C0",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"02",X"01",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"02",X"02",X"00",X"5B",X"A0",X"60",X"B8",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"07",X"06",X"00",X"5B",X"F0",X"50",X"18",X"20",X"28",X"60",X"D0",X"60",X"28",X"18",X"A8",X"61",
		X"05",X"00",X"A0",X"5B",X"F0",X"50",X"C0",X"30",X"E0",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"04",X"00",X"C0",X"5B",X"F0",X"50",X"C0",X"30",X"E0",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"04",X"00",X"E0",X"5B",X"F0",X"50",X"E0",X"30",X"C8",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"03",X"01",X"40",X"5B",X"F0",X"50",X"E0",X"30",X"C8",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"48",X"10",X"40",X"DF",X"3F",
		X"04",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"28",X"40",X"E8",X"3F",
		X"0E",X"00",X"A0",X"5B",X"08",X"30",X"18",X"30",X"38",X"40",X"EC",X"30",X"D4",X"2E",X"CB",X"20",
		X"04",X"02",X"80",X"5B",X"00",X"60",X"18",X"50",X"38",X"50",X"F4",X"08",X"DC",X"5E",X"A1",X"5C",
		X"04",X"06",X"00",X"5B",X"08",X"00",X"28",X"40",X"38",X"40",X"04",X"60",X"F0",X"66",X"A1",X"5A",
		X"03",X"06",X"00",X"5B",X"28",X"40",X"38",X"40",X"08",X"00",X"04",X"50",X"F4",X"62",X"A4",X"57",
		X"03",X"06",X"00",X"5B",X"08",X"10",X"28",X"50",X"38",X"40",X"04",X"48",X"F4",X"64",X"9A",X"62",
		X"03",X"06",X"00",X"5B",X"08",X"20",X"28",X"50",X"38",X"40",X"04",X"38",X"F8",X"60",X"96",X"66",
		X"05",X"04",X"00",X"5B",X"08",X"30",X"28",X"50",X"38",X"50",X"FC",X"20",X"F8",X"62",X"92",X"6E",
		X"04",X"01",X"40",X"5B",X"08",X"40",X"28",X"40",X"38",X"40",X"F8",X"60",X"F4",X"0C",X"90",X"71",
		X"03",X"03",X"00",X"5B",X"A0",X"70",X"E8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"01",X"03",X"00",X"5B",X"A0",X"70",X"F0",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"A0",X"70",X"F0",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"01",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"F8",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"06",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"01",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"07",X"00",X"A0",X"5B",X"90",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"02",X"00",X"70",X"5B",X"90",X"70",X"F8",X"60",X"F8",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"04",X"02",X"80",X"5B",X"90",X"70",X"E0",X"70",X"00",X"60",X"10",X"10",X"1C",X"56",X"3A",X"49",
		X"02",X"02",X"00",X"5B",X"98",X"70",X"E0",X"70",X"00",X"60",X"10",X"10",X"1C",X"56",X"3A",X"49",
		X"04",X"05",X"00",X"5B",X"98",X"60",X"F0",X"60",X"D8",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C",
		X"02",X"05",X"00",X"5B",X"D0",X"60",X"F0",X"60",X"A0",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C",
		X"03",X"04",X"00",X"5B",X"F0",X"60",X"C8",X"60",X"A0",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C",
		X"09",X"04",X"00",X"5B",X"20",X"50",X"18",X"20",X"40",X"30",X"F8",X"60",X"C0",X"60",X"B2",X"5A",
		X"04",X"05",X"00",X"5B",X"C8",X"60",X"B8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41",
		X"02",X"05",X"00",X"5B",X"C8",X"60",X"B8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41",
		X"03",X"05",X"00",X"5B",X"B8",X"60",X"C8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41",
		X"03",X"01",X"C0",X"5B",X"10",X"50",X"28",X"40",X"30",X"30",X"08",X"30",X"F0",X"64",X"8E",X"70",
		X"03",X"01",X"80",X"5B",X"10",X"50",X"28",X"50",X"38",X"30",X"04",X"28",X"F4",X"5E",X"8C",X"76",
		X"04",X"02",X"80",X"5B",X"08",X"30",X"28",X"40",X"30",X"20",X"08",X"40",X"F4",X"5C",X"90",X"70",
		X"02",X"04",X"00",X"5B",X"10",X"30",X"20",X"50",X"38",X"40",X"00",X"38",X"F0",X"5A",X"95",X"69",
		X"02",X"07",X"00",X"5B",X"20",X"40",X"28",X"40",X"18",X"10",X"00",X"48",X"F0",X"60",X"98",X"69",
		X"02",X"06",X"00",X"5B",X"18",X"30",X"28",X"40",X"20",X"10",X"00",X"48",X"F0",X"5E",X"9C",X"68",
		X"0A",X"03",X"00",X"5B",X"F8",X"40",X"20",X"50",X"30",X"50",X"F0",X"20",X"DC",X"4C",X"AE",X"66",
		X"07",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"28",X"08",X"4E",X"EB",X"0C",
		X"07",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"38",X"0C",X"3E",X"F1",X"1A",
		X"02",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"E8",X"F2",X"03",X"3F",
		X"03",X"00",X"04",X"5B",X"F8",X"30",X"18",X"40",X"40",X"30",X"E4",X"20",X"18",X"04",X"88",X"76",
		X"01",X"03",X"00",X"5B",X"20",X"50",X"18",X"10",X"30",X"40",X"F8",X"78",X"E0",X"74",X"98",X"6C",
		X"16",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"24",X"E5",X"3B",
		X"09",X"02",X"80",X"5B",X"F8",X"70",X"20",X"50",X"28",X"50",X"C0",X"68",X"18",X"06",X"A4",X"5E",
		X"09",X"02",X"80",X"5B",X"F0",X"60",X"18",X"60",X"20",X"40",X"D8",X"60",X"20",X"0C",X"9D",X"61",
		X"05",X"03",X"00",X"5B",X"18",X"50",X"20",X"50",X"38",X"30",X"F0",X"60",X"D0",X"66",X"A6",X"53",
		X"08",X"02",X"00",X"5B",X"18",X"60",X"28",X"50",X"40",X"40",X"F0",X"60",X"C8",X"62",X"9D",X"61",
		X"09",X"01",X"C0",X"5B",X"B8",X"60",X"D0",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"06",X"01",X"00",X"5B",X"B0",X"60",X"C8",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"04",X"00",X"A0",X"5B",X"B0",X"60",X"C0",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"05",X"00",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"08",X"00",X"28",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"09",X"00",X"18",X"5B",X"00",X"40",X"20",X"30",X"38",X"30",X"E4",X"28",X"08",X"F8",X"91",X"65",
		X"01",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"20",X"14",X"30",X"E6",X"27",
		X"05",X"08",X"00",X"5B",X"20",X"60",X"28",X"30",X"40",X"30",X"FC",X"58",X"E4",X"70",X"A7",X"4B",
		X"07",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"40",X"F4",X"4C",X"E7",X"23",
		X"05",X"01",X"80",X"5B",X"F8",X"70",X"30",X"60",X"30",X"30",X"E8",X"60",X"08",X"FC",X"AC",X"48",
		X"07",X"00",X"20",X"5B",X"08",X"30",X"28",X"50",X"50",X"40",X"F0",X"48",X"C8",X"68",X"A8",X"47",
		X"07",X"00",X"E0",X"5B",X"10",X"40",X"28",X"40",X"50",X"50",X"F0",X"40",X"D0",X"1A",X"DE",X"3A",
		X"02",X"01",X"40",X"5B",X"F0",X"60",X"18",X"40",X"20",X"40",X"D0",X"68",X"2C",X"18",X"C7",X"25",
		X"03",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"30",X"FC",X"F0",X"FB",X"41",
		X"03",X"07",X"00",X"5B",X"10",X"40",X"20",X"60",X"38",X"30",X"F8",X"30",X"F4",X"5E",X"A1",X"5C",
		X"04",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"10",X"20",X"4E",X"FA",X"53",
		X"0A",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"18",X"44",X"FC",X"5A",
		X"06",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"14",X"40",X"FB",X"5D",
		X"08",X"01",X"40",X"5B",X"C0",X"30",X"E0",X"40",X"F8",X"60",X"14",X"58",X"24",X"48",X"00",X"00",
		X"0C",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"42",X"FE",X"3F",
		X"02",X"00",X"38",X"5B",X"08",X"40",X"20",X"30",X"38",X"30",X"DC",X"48",X"BC",X"58",X"A4",X"54",
		X"04",X"00",X"60",X"5B",X"D0",X"60",X"10",X"70",X"20",X"30",X"BC",X"60",X"1C",X"08",X"A1",X"5D",
		X"04",X"00",X"A0",X"5B",X"D0",X"50",X"10",X"60",X"18",X"50",X"BC",X"60",X"20",X"0E",X"A3",X"5C",
		X"13",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"04",X"28",X"E3",X"27",
		X"14",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"30",X"04",X"12",X"DE",X"56",
		X"01",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"28",X"F4",X"1E",X"DC",X"49",
		X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"0C",X"62",X"E2",X"37",
		X"01",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"20",X"10",X"36",X"F9",X"44",
		X"0A",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"28",X"0C",X"44",X"E7",X"1B",
		X"07",X"04",X"00",X"5B",X"20",X"50",X"40",X"60",X"58",X"50",X"00",X"58",X"DC",X"54",X"A7",X"4D",
		X"0A",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"58",X"EC",X"00",X"21",X"30",
		X"05",X"05",X"00",X"5B",X"20",X"50",X"40",X"50",X"48",X"40",X"00",X"40",X"DC",X"60",X"B9",X"37",
		X"04",X"03",X"80",X"5B",X"D8",X"40",X"B8",X"40",X"F8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"03",X"02",X"00",X"5B",X"F0",X"40",X"B0",X"40",X"D8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"05",X"01",X"C0",X"5B",X"B0",X"40",X"F0",X"40",X"D8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"07",X"01",X"40",X"5B",X"F0",X"40",X"B0",X"40",X"D0",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"04",X"00",X"C0",X"5B",X"98",X"60",X"C8",X"60",X"08",X"40",X"18",X"30",X"28",X"44",X"2E",X"25",
		X"04",X"02",X"80",X"5B",X"A0",X"60",X"C8",X"60",X"08",X"40",X"18",X"30",X"28",X"44",X"2E",X"25",
		X"04",X"02",X"00",X"5B",X"A0",X"60",X"C0",X"60",X"00",X"40",X"18",X"30",X"28",X"44",X"2E",X"25",
		X"04",X"00",X"10",X"5B",X"A0",X"60",X"B0",X"50",X"20",X"40",X"F8",X"18",X"1C",X"52",X"00",X"00",
		X"03",X"00",X"14",X"5B",X"A0",X"60",X"B0",X"50",X"18",X"40",X"F8",X"18",X"1C",X"52",X"00",X"00",
		X"05",X"00",X"1C",X"5B",X"A0",X"60",X"B0",X"50",X"20",X"40",X"F8",X"18",X"1C",X"52",X"00",X"00",
		X"04",X"00",X"28",X"5B",X"A0",X"60",X"B0",X"50",X"18",X"40",X"F8",X"18",X"1C",X"52",X"00",X"00",
		X"04",X"02",X"80",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"02",X"80",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"03",X"01",X"C0",X"5B",X"A0",X"60",X"E8",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"02",X"80",X"5B",X"A0",X"60",X"E0",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"03",X"00",X"5B",X"A8",X"60",X"E0",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"03",X"02",X"80",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"03",X"02",X"00",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"01",X"C0",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"00",X"E0",X"5B",X"A8",X"60",X"D0",X"60",X"E0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"00",X"80",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"00",X"C0",X"5B",X"A8",X"60",X"D0",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"00",X"70",X"5B",X"A8",X"60",X"D0",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"00",X"50",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"07",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"FC",X"1C",X"D2",X"28",
		X"0C",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"38",X"04",X"18",X"B4",X"55",
		X"02",X"00",X"C0",X"5B",X"F8",X"40",X"30",X"70",X"20",X"20",X"C4",X"38",X"10",X"FC",X"A3",X"5D",
		X"02",X"01",X"40",X"5B",X"F8",X"60",X"28",X"50",X"28",X"50",X"B0",X"68",X"1C",X"06",X"A3",X"58",
		X"03",X"01",X"C0",X"5B",X"10",X"50",X"28",X"40",X"30",X"30",X"08",X"30",X"F0",X"64",X"8E",X"70",
		X"03",X"01",X"80",X"5B",X"10",X"50",X"28",X"50",X"38",X"30",X"04",X"28",X"F4",X"5E",X"8C",X"76",
		X"04",X"02",X"80",X"5B",X"08",X"30",X"28",X"40",X"30",X"20",X"08",X"40",X"F4",X"5C",X"90",X"70",
		X"02",X"04",X"00",X"5B",X"10",X"30",X"20",X"50",X"38",X"40",X"00",X"38",X"F0",X"5A",X"95",X"69",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"08",X"4E",X"E4",X"19",
		X"0E",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"50",X"10",X"66",X"F6",X"49",
		X"01",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"30",X"20",X"E4",X"60",X"CC",X"68",X"A5",X"5F",
		X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"28",X"10",X"E4",X"58",X"D0",X"60",X"A5",X"5F",
		X"01",X"02",X"80",X"5B",X"E0",X"60",X"18",X"40",X"20",X"40",X"D0",X"60",X"24",X"12",X"A8",X"5B",
		X"01",X"02",X"00",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"20",X"0A",X"A3",X"63",
		X"01",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D0",X"68",X"20",X"0A",X"A5",X"61",
		X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"24",X"12",X"A2",X"69",
		X"01",X"01",X"40",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D4",X"68",X"1C",X"0A",X"A0",X"6E",
		X"02",X"00",X"E0",X"5B",X"18",X"60",X"20",X"20",X"20",X"10",X"E0",X"60",X"D4",X"68",X"A0",X"6E",
		X"01",X"00",X"E0",X"5B",X"18",X"60",X"18",X"20",X"30",X"20",X"E4",X"60",X"D4",X"6A",X"A3",X"63",
		X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"30",X"20",X"E4",X"60",X"CC",X"68",X"A5",X"5F",
		X"03",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"28",X"10",X"E4",X"58",X"D0",X"60",X"A5",X"5F",
		X"01",X"02",X"00",X"5B",X"E0",X"60",X"18",X"40",X"28",X"40",X"D0",X"60",X"24",X"10",X"A9",X"59",
		X"03",X"02",X"00",X"5B",X"E0",X"60",X"18",X"40",X"20",X"40",X"D0",X"60",X"24",X"12",X"A8",X"5B",
		X"01",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"20",X"0A",X"A3",X"63",
		X"03",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D0",X"68",X"20",X"0A",X"A5",X"61",
		X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"24",X"12",X"A2",X"69",
		X"04",X"01",X"40",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D4",X"68",X"1C",X"0A",X"A0",X"6E",
		X"03",X"00",X"C0",X"5B",X"18",X"60",X"20",X"20",X"20",X"10",X"E0",X"60",X"D4",X"68",X"A0",X"6E",
		X"04",X"00",X"E0",X"5B",X"18",X"60",X"18",X"20",X"30",X"20",X"E4",X"60",X"D4",X"6A",X"A3",X"63",
		X"03",X"02",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"02",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"02",X"00",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"02",X"01",X"C0",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"05",X"00",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"02",X"00",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"06",X"00",X"70",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"13",X"00",X"A0",X"5B",X"08",X"30",X"18",X"30",X"38",X"40",X"EC",X"30",X"D4",X"2E",X"CB",X"20",
		X"04",X"02",X"80",X"5B",X"00",X"60",X"18",X"50",X"38",X"50",X"F4",X"08",X"DC",X"5E",X"A1",X"5C",
		X"0B",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"40",X"20",X"38",X"E3",X"29",
		X"04",X"00",X"A0",X"5B",X"00",X"30",X"18",X"20",X"38",X"40",X"FC",X"60",X"E0",X"2A",X"A1",X"54",
		X"03",X"00",X"C0",X"5B",X"08",X"30",X"20",X"30",X"20",X"10",X"FC",X"68",X"E8",X"1C",X"A2",X"50",
		X"02",X"00",X"C0",X"5B",X"08",X"30",X"20",X"40",X"20",X"10",X"FC",X"68",X"E0",X"24",X"9B",X"5B",
		X"04",X"06",X"00",X"5B",X"10",X"40",X"18",X"40",X"30",X"30",X"F8",X"68",X"DC",X"62",X"A8",X"50",
		X"01",X"06",X"00",X"5B",X"10",X"20",X"18",X"40",X"30",X"40",X"F8",X"68",X"D4",X"6E",X"AC",X"55",
		X"03",X"06",X"00",X"5B",X"20",X"50",X"18",X"10",X"30",X"40",X"F8",X"70",X"D0",X"6A",X"AC",X"58",
		X"12",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"00",X"1E",X"C1",X"48",
		X"02",X"00",X"C0",X"5B",X"F8",X"50",X"20",X"60",X"40",X"60",X"C4",X"48",X"EC",X"FE",X"BA",X"43",
		X"02",X"00",X"A0",X"5B",X"F8",X"40",X"18",X"60",X"40",X"60",X"C0",X"68",X"E8",X"00",X"A9",X"5E",
		X"02",X"00",X"60",X"5B",X"A0",X"60",X"A8",X"60",X"F8",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"02",X"00",X"40",X"5B",X"A0",X"60",X"A8",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"02",X"00",X"50",X"5B",X"A0",X"60",X"A8",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"05",X"00",X"E0",X"5B",X"A0",X"60",X"B0",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"04",X"01",X"40",X"5B",X"A0",X"60",X"C0",X"60",X"E8",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"06",X"01",X"C0",X"5B",X"A8",X"60",X"C8",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"03",X"01",X"C0",X"5B",X"A8",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"03",X"00",X"E0",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"02",X"00",X"60",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"02",X"01",X"00",X"5B",X"18",X"60",X"28",X"40",X"10",X"00",X"F0",X"48",X"BC",X"64",X"AC",X"59",
		X"02",X"01",X"40",X"5B",X"10",X"60",X"20",X"40",X"18",X"10",X"F0",X"48",X"BC",X"62",X"AF",X"56",
		X"02",X"01",X"80",X"5B",X"10",X"50",X"20",X"30",X"20",X"10",X"EC",X"48",X"C0",X"5E",X"B0",X"56",
		X"03",X"01",X"40",X"5B",X"F0",X"50",X"10",X"60",X"20",X"50",X"C0",X"60",X"10",X"02",X"B6",X"51",
		X"02",X"01",X"40",X"5B",X"E8",X"60",X"18",X"60",X"28",X"50",X"C4",X"60",X"04",X"00",X"B8",X"4A",
		X"04",X"01",X"40",X"5B",X"18",X"60",X"10",X"00",X"20",X"30",X"E8",X"58",X"C8",X"62",X"B5",X"54",
		X"03",X"00",X"E0",X"5B",X"00",X"00",X"18",X"60",X"30",X"50",X"E4",X"60",X"CC",X"58",X"B5",X"56",
		X"04",X"00",X"C0",X"5B",X"00",X"00",X"18",X"60",X"28",X"40",X"E4",X"60",X"D0",X"5C",X"B2",X"59",
		X"03",X"00",X"80",X"5B",X"E8",X"60",X"10",X"60",X"20",X"20",X"CC",X"60",X"04",X"FC",X"B2",X"55",
		X"03",X"03",X"80",X"5B",X"90",X"70",X"F0",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"04",X"00",X"5B",X"90",X"70",X"F8",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"05",X"00",X"5B",X"90",X"70",X"F8",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"02",X"80",X"5B",X"90",X"70",X"F0",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"02",X"80",X"5B",X"98",X"70",X"E8",X"50",X"F8",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"05",X"01",X"80",X"5B",X"A0",X"70",X"E0",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"05",X"01",X"80",X"5B",X"A0",X"70",X"D8",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"06",X"01",X"40",X"5B",X"A0",X"70",X"D8",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"C0",X"5B",X"08",X"40",X"20",X"40",X"38",X"50",X"E4",X"48",X"DC",X"44",X"BD",X"3D",
		X"06",X"03",X"00",X"5B",X"18",X"40",X"28",X"50",X"20",X"20",X"FC",X"68",X"C4",X"60",X"A3",X"64",
		X"03",X"01",X"80",X"5B",X"10",X"10",X"28",X"60",X"38",X"40",X"FC",X"60",X"C0",X"62",X"A3",X"60",
		X"08",X"01",X"00",X"5B",X"28",X"60",X"18",X"10",X"30",X"30",X"00",X"60",X"C0",X"60",X"A0",X"68",
		X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"20",X"FC",X"20",X"DE",X"48",
		X"02",X"04",X"00",X"5B",X"20",X"50",X"30",X"40",X"18",X"10",X"F8",X"68",X"E0",X"6C",X"98",X"6C",
		X"04",X"07",X"00",X"3D",X"08",X"30",X"10",X"20",X"38",X"50",X"F0",X"48",X"E4",X"1C",X"A9",X"63",
		X"03",X"06",X"00",X"38",X"10",X"40",X"18",X"20",X"38",X"50",X"F0",X"50",X"D8",X"22",X"A9",X"5D",
		X"04",X"06",X"00",X"2F",X"10",X"20",X"18",X"30",X"40",X"60",X"F0",X"48",X"DC",X"1A",X"AC",X"5F",
		X"04",X"06",X"00",X"2C",X"00",X"10",X"18",X"50",X"40",X"60",X"EC",X"50",X"B0",X"56",X"E5",X"0D",
		X"04",X"07",X"00",X"2A",X"10",X"20",X"18",X"60",X"38",X"50",X"E8",X"58",X"DC",X"1A",X"B9",X"44",
		X"05",X"02",X"00",X"2C",X"08",X"40",X"20",X"40",X"38",X"50",X"E0",X"60",X"E4",X"0C",X"AF",X"42",
		X"04",X"04",X"00",X"2A",X"08",X"40",X"10",X"30",X"30",X"40",X"E0",X"68",X"E4",X"02",X"B1",X"54",
		X"06",X"06",X"00",X"2B",X"08",X"50",X"18",X"40",X"38",X"40",X"E0",X"60",X"E0",X"08",X"B3",X"54",
		X"05",X"06",X"00",X"2D",X"08",X"50",X"20",X"50",X"38",X"40",X"DC",X"60",X"DC",X"10",X"B1",X"53",
		X"04",X"03",X"80",X"34",X"00",X"20",X"18",X"30",X"30",X"50",X"DC",X"48",X"E4",X"0A",X"B4",X"43",
		X"06",X"01",X"C0",X"41",X"F8",X"60",X"20",X"60",X"38",X"60",X"F8",X"08",X"D8",X"5C",X"A3",X"50",
		X"04",X"01",X"00",X"62",X"18",X"60",X"10",X"10",X"38",X"70",X"F4",X"70",X"D4",X"5A",X"9C",X"5A",
		X"03",X"03",X"80",X"6E",X"00",X"60",X"18",X"60",X"38",X"50",X"E4",X"60",X"F0",X"04",X"AA",X"50",
		X"02",X"02",X"80",X"6F",X"00",X"50",X"20",X"50",X"30",X"40",X"EC",X"60",X"EC",X"00",X"AC",X"4E",
		X"03",X"01",X"C0",X"67",X"08",X"50",X"20",X"50",X"40",X"50",X"F0",X"58",X"E8",X"06",X"A7",X"57",
		X"02",X"01",X"40",X"81",X"08",X"50",X"20",X"40",X"40",X"60",X"F4",X"68",X"EC",X"0A",X"9F",X"60",
		X"03",X"00",X"E0",X"83",X"08",X"60",X"28",X"50",X"40",X"60",X"F8",X"70",X"E8",X"0A",X"9D",X"60",
		X"02",X"00",X"E0",X"88",X"08",X"40",X"20",X"40",X"40",X"60",X"F8",X"58",X"F0",X"0C",X"92",X"73",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"03",X"00",X"47",X"00",X"00",X"20",X"60",X"38",X"70",X"04",X"60",X"BC",X"6E",X"A5",X"76",
		X"04",X"04",X"00",X"45",X"00",X"60",X"20",X"60",X"40",X"70",X"FC",X"08",X"BC",X"68",X"AA",X"65",
		X"04",X"03",X"80",X"3F",X"00",X"00",X"20",X"60",X"40",X"70",X"00",X"60",X"BC",X"68",X"A6",X"75",
		X"06",X"05",X"00",X"39",X"00",X"00",X"20",X"60",X"40",X"70",X"00",X"60",X"C0",X"5A",X"AB",X"67",
		X"05",X"03",X"80",X"38",X"00",X"50",X"20",X"60",X"40",X"60",X"FC",X"00",X"BC",X"62",X"AD",X"60",
		X"05",X"02",X"00",X"35",X"F8",X"60",X"20",X"60",X"40",X"60",X"F4",X"00",X"BC",X"62",X"AC",X"60",
		X"06",X"01",X"C0",X"31",X"00",X"60",X"20",X"60",X"48",X"60",X"F8",X"00",X"BC",X"5E",X"A8",X"66",
		X"05",X"01",X"80",X"31",X"00",X"60",X"20",X"60",X"40",X"50",X"F4",X"00",X"BC",X"58",X"AB",X"5A",
		X"05",X"01",X"40",X"33",X"08",X"60",X"20",X"50",X"40",X"40",X"C0",X"58",X"F0",X"06",X"A9",X"57",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"40",X"14",X"3C",X"BE",X"6C",
		X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"50",X"0C",X"28",X"CB",X"44",
		X"04",X"02",X"00",X"4B",X"10",X"30",X"28",X"60",X"38",X"60",X"F4",X"48",X"C4",X"56",X"A3",X"59",
		X"04",X"05",X"00",X"57",X"08",X"10",X"20",X"50",X"30",X"50",X"F4",X"50",X"E0",X"66",X"9B",X"70",
		X"04",X"05",X"00",X"5D",X"10",X"20",X"18",X"50",X"30",X"50",X"F0",X"48",X"E4",X"58",X"97",X"74",
		X"04",X"05",X"00",X"61",X"18",X"50",X"18",X"20",X"30",X"60",X"F0",X"50",X"E8",X"5C",X"95",X"75",
		X"03",X"05",X"00",X"63",X"18",X"50",X"18",X"20",X"30",X"50",X"F0",X"60",X"E4",X"5E",X"97",X"72",
		X"04",X"05",X"00",X"65",X"18",X"40",X"20",X"40",X"38",X"50",X"EC",X"60",X"E0",X"6A",X"9B",X"6D",
		X"03",X"03",X"80",X"67",X"20",X"60",X"30",X"50",X"18",X"10",X"E8",X"58",X"DC",X"60",X"9F",X"6E",
		X"03",X"03",X"80",X"64",X"20",X"50",X"10",X"10",X"30",X"50",X"E8",X"58",X"DC",X"64",X"A0",X"6C",
		X"03",X"02",X"00",X"61",X"08",X"10",X"20",X"50",X"40",X"60",X"E8",X"50",X"DC",X"58",X"A3",X"62",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"40",X"08",X"4A",X"C9",X"48",
		X"05",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"E0",X"10",X"01",X"19",
		X"04",X"01",X"00",X"35",X"08",X"50",X"28",X"70",X"40",X"70",X"F0",X"08",X"C0",X"70",X"9B",X"68",
		X"03",X"02",X"00",X"31",X"10",X"70",X"20",X"50",X"38",X"70",X"04",X"10",X"C0",X"74",X"99",X"6B",
		X"04",X"05",X"00",X"31",X"10",X"60",X"28",X"60",X"38",X"70",X"E0",X"48",X"E0",X"28",X"9F",X"67",
		X"04",X"06",X"00",X"32",X"08",X"60",X"28",X"40",X"38",X"50",X"E0",X"70",X"E4",X"18",X"A0",X"64",
		X"06",X"06",X"00",X"38",X"00",X"60",X"28",X"40",X"38",X"60",X"F0",X"58",X"E8",X"18",X"9A",X"67",
		X"02",X"05",X"00",X"47",X"00",X"50",X"20",X"30",X"38",X"60",X"F8",X"58",X"F0",X"0A",X"96",X"69",
		X"04",X"03",X"80",X"60",X"00",X"50",X"20",X"50",X"38",X"60",X"F8",X"58",X"F4",X"0A",X"94",X"6B",
		X"02",X"01",X"C0",X"7A",X"08",X"50",X"20",X"50",X"38",X"60",X"F8",X"58",X"EC",X"04",X"91",X"70",
		X"03",X"01",X"C0",X"8E",X"00",X"50",X"20",X"60",X"40",X"60",X"F8",X"60",X"F4",X"0C",X"91",X"6D",
		X"02",X"01",X"40",X"93",X"00",X"50",X"20",X"50",X"40",X"60",X"F4",X"58",X"F4",X"08",X"8E",X"77",
		X"02",X"00",X"C0",X"94",X"00",X"60",X"20",X"30",X"40",X"60",X"EC",X"58",X"F0",X"06",X"90",X"73",
		X"03",X"00",X"C0",X"9D",X"00",X"60",X"38",X"60",X"30",X"40",X"E4",X"68",X"F8",X"FA",X"96",X"69",
		X"06",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"60",X"10",X"FC",X"E7",X"24",
		X"04",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"38",X"24",X"3A",X"E2",X"30",
		X"07",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"48",X"1C",X"16",X"DF",X"2F",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"C0",X"5B",X"08",X"50",X"20",X"60",X"38",X"60",X"F4",X"58",X"F4",X"18",X"8C",X"7F",
		X"03",X"07",X"00",X"4A",X"00",X"40",X"20",X"50",X"38",X"50",X"F8",X"18",X"F0",X"58",X"95",X"78",
		X"05",X"06",X"00",X"4C",X"00",X"40",X"20",X"40",X"38",X"50",X"F8",X"10",X"EC",X"52",X"A1",X"68",
		X"04",X"06",X"00",X"42",X"00",X"50",X"18",X"40",X"38",X"50",X"E8",X"50",X"F0",X"10",X"A4",X"74",
		X"05",X"06",X"00",X"3B",X"00",X"50",X"18",X"30",X"40",X"60",X"F4",X"10",X"E8",X"58",X"A8",X"73",
		X"04",X"06",X"00",X"3A",X"00",X"50",X"18",X"20",X"40",X"60",X"E8",X"58",X"F4",X"0C",X"A9",X"6D",
		X"04",X"07",X"00",X"39",X"00",X"50",X"20",X"20",X"40",X"60",X"E8",X"50",X"E8",X"16",X"A8",X"60",
		X"03",X"03",X"80",X"3D",X"00",X"50",X"20",X"20",X"40",X"60",X"E4",X"60",X"E8",X"0C",X"B5",X"44",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"40",X"F0",X"24",X"DB",X"23",
		X"2A",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"01",X"80",X"5C",X"00",X"00",X"10",X"50",X"30",X"70",X"04",X"68",X"BC",X"6A",X"A5",X"6E",
		X"04",X"02",X"80",X"58",X"10",X"60",X"08",X"00",X"28",X"70",X"04",X"70",X"B8",X"72",X"A5",X"6D",
		X"04",X"03",X"00",X"55",X"08",X"70",X"10",X"50",X"28",X"60",X"B8",X"70",X"0C",X"02",X"A5",X"6F",
		X"03",X"03",X"00",X"55",X"10",X"60",X"08",X"00",X"28",X"60",X"04",X"68",X"B8",X"6C",X"A7",X"6E",
		X"04",X"03",X"80",X"5A",X"10",X"50",X"28",X"60",X"08",X"00",X"04",X"68",X"BC",X"66",X"A7",X"70",
		X"04",X"04",X"00",X"5D",X"08",X"70",X"10",X"50",X"28",X"60",X"BC",X"70",X"0C",X"02",X"A7",X"6E",
		X"03",X"03",X"00",X"63",X"10",X"50",X"28",X"60",X"08",X"00",X"04",X"70",X"C0",X"5C",X"A7",X"74",
		X"04",X"03",X"00",X"68",X"00",X"60",X"10",X"50",X"28",X"60",X"BC",X"70",X"0C",X"02",X"AC",X"65",
		X"03",X"02",X"80",X"72",X"08",X"40",X"08",X"00",X"28",X"40",X"04",X"58",X"C0",X"6E",X"AD",X"68",
		X"02",X"01",X"00",X"7A",X"00",X"60",X"18",X"30",X"30",X"40",X"C0",X"78",X"F0",X"04",X"AD",X"6F",
		X"03",X"00",X"C0",X"7F",X"00",X"60",X"18",X"20",X"38",X"70",X"C0",X"70",X"F4",X"FC",X"AF",X"66",
		X"02",X"00",X"C0",X"88",X"00",X"50",X"28",X"50",X"30",X"50",X"F0",X"08",X"C4",X"62",X"AC",X"6D",
		X"04",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"58",X"E4",X"1C",X"C4",X"4F",
		X"06",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"40",X"F8",X"24",X"C9",X"25",
		X"08",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"38",X"04",X"1E",X"DC",X"3D",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"03",X"80",X"4B",X"18",X"60",X"18",X"10",X"30",X"50",X"08",X"60",X"B4",X"60",X"A0",X"6C",
		X"05",X"02",X"80",X"44",X"20",X"70",X"30",X"60",X"10",X"00",X"08",X"60",X"B0",X"62",X"99",X"71",
		X"04",X"01",X"80",X"41",X"08",X"60",X"20",X"70",X"38",X"50",X"A8",X"68",X"04",X"00",X"A1",X"5B",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"48",X"F0",X"2A",X"CC",X"2D",
		X"04",X"03",X"80",X"33",X"00",X"50",X"20",X"60",X"38",X"70",X"F0",X"10",X"DC",X"6C",X"96",X"75",
		X"04",X"03",X"80",X"33",X"00",X"60",X"28",X"60",X"38",X"70",X"F4",X"08",X"DC",X"72",X"98",X"6F",
		X"04",X"02",X"00",X"33",X"00",X"60",X"28",X"60",X"38",X"60",X"DC",X"68",X"9C",X"60",X"F5",X"02",
		X"11",X"00",X"E0",X"35",X"00",X"50",X"20",X"30",X"40",X"70",X"F4",X"28",X"D0",X"58",X"9F",X"58",
		X"07",X"01",X"80",X"34",X"00",X"50",X"28",X"50",X"38",X"60",X"F4",X"38",X"D0",X"42",X"A1",X"56",
		X"09",X"01",X"40",X"34",X"08",X"60",X"30",X"50",X"40",X"60",X"F0",X"38",X"D4",X"30",X"A3",X"52",
		X"16",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"38",X"F8",X"20",X"C9",X"36",
		X"03",X"07",X"00",X"46",X"08",X"10",X"20",X"60",X"28",X"50",X"00",X"60",X"BC",X"6E",X"A5",X"6D",
		X"05",X"06",X"00",X"45",X"00",X"60",X"20",X"60",X"28",X"60",X"00",X"08",X"C4",X"60",X"AC",X"68",
		X"03",X"06",X"00",X"4A",X"00",X"60",X"20",X"50",X"28",X"60",X"F4",X"10",X"C8",X"5C",X"B3",X"67",
		X"04",X"06",X"00",X"4C",X"00",X"60",X"20",X"50",X"28",X"60",X"F0",X"10",X"CC",X"62",X"B6",X"61",
		X"03",X"07",X"00",X"55",X"F8",X"50",X"20",X"50",X"30",X"50",X"F4",X"10",X"D8",X"60",X"B0",X"6C",
		X"04",X"05",X"00",X"67",X"00",X"00",X"18",X"50",X"28",X"40",X"F8",X"50",X"E4",X"58",X"A7",X"67",
		X"03",X"05",X"00",X"75",X"10",X"50",X"20",X"40",X"30",X"40",X"F4",X"48",X"E4",X"60",X"9E",X"6F",
		X"03",X"02",X"80",X"79",X"08",X"20",X"18",X"50",X"38",X"50",X"EC",X"50",X"E4",X"5E",X"9E",X"6A",
		X"03",X"01",X"C0",X"7C",X"08",X"10",X"10",X"50",X"38",X"50",X"E8",X"60",X"DC",X"68",X"A0",X"6D",
		X"04",X"01",X"C0",X"81",X"10",X"50",X"10",X"10",X"40",X"60",X"E4",X"68",X"D4",X"68",X"A2",X"70",
		X"03",X"01",X"C0",X"86",X"10",X"20",X"10",X"40",X"38",X"60",X"E4",X"60",X"D4",X"66",X"A2",X"71",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"A0",X"56",X"08",X"60",X"20",X"70",X"28",X"40",X"AC",X"78",X"0C",X"FC",X"9A",X"6C",
		X"03",X"03",X"80",X"47",X"08",X"10",X"20",X"60",X"38",X"60",X"04",X"58",X"BC",X"6E",X"A4",X"75",
		X"04",X"07",X"00",X"3E",X"08",X"00",X"20",X"60",X"40",X"70",X"FC",X"60",X"C8",X"74",X"A8",X"73",
		X"03",X"06",X"00",X"38",X"F8",X"50",X"20",X"50",X"40",X"60",X"D8",X"60",X"F8",X"00",X"AC",X"64",
		X"03",X"06",X"00",X"35",X"00",X"50",X"20",X"40",X"40",X"50",X"F0",X"10",X"E0",X"5E",X"A8",X"5E",
		X"02",X"02",X"00",X"5A",X"F8",X"30",X"20",X"50",X"38",X"50",X"E0",X"58",X"08",X"FC",X"A9",X"4C",
		X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"40",X"14",X"40",X"E9",X"24",
		X"05",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"50",X"14",X"42",X"EE",X"19",
		X"03",X"02",X"80",X"4C",X"08",X"50",X"20",X"50",X"40",X"40",X"EC",X"50",X"EC",X"0E",X"A3",X"5C",
		X"02",X"05",X"00",X"2F",X"00",X"50",X"18",X"60",X"40",X"50",X"EC",X"58",X"EC",X"0E",X"A5",X"5F",
		X"05",X"05",X"00",X"2E",X"00",X"50",X"20",X"50",X"40",X"50",X"E8",X"48",X"E4",X"16",X"AB",X"5A",
		X"05",X"04",X"00",X"2D",X"00",X"40",X"20",X"50",X"40",X"50",X"E4",X"48",X"E8",X"1C",X"AF",X"62",
		X"06",X"03",X"80",X"2D",X"F8",X"50",X"20",X"40",X"40",X"50",X"DC",X"50",X"F0",X"0A",X"BA",X"5D",
		X"05",X"03",X"00",X"30",X"F8",X"40",X"20",X"40",X"40",X"50",X"DC",X"50",X"F0",X"04",X"BB",X"67",
		X"05",X"02",X"80",X"30",X"F8",X"50",X"20",X"50",X"40",X"50",X"F4",X"08",X"D0",X"5E",X"B7",X"65",
		X"05",X"03",X"80",X"38",X"F8",X"50",X"20",X"50",X"40",X"60",X"F8",X"08",X"CC",X"5C",X"B3",X"64",
		X"03",X"02",X"80",X"55",X"F8",X"60",X"20",X"60",X"40",X"60",X"C8",X"60",X"B0",X"60",X"F8",X"01",
		X"03",X"00",X"E0",X"69",X"00",X"50",X"20",X"60",X"40",X"50",X"C4",X"60",X"F0",X"02",X"AA",X"64",
		X"02",X"00",X"70",X"77",X"00",X"40",X"20",X"50",X"38",X"40",X"C0",X"68",X"F8",X"FE",X"A7",X"5F",
		X"02",X"00",X"80",X"85",X"F8",X"60",X"18",X"60",X"38",X"50",X"C4",X"68",X"0C",X"FE",X"A3",X"62",
		X"0E",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"10",X"14",X"14",X"BC",X"41",
		X"01",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"F8",X"1C",X"DF",X"13",
		X"02",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"F4",X"28",X"E7",X"11",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"C0",X"3C",X"F0",X"60",X"18",X"60",X"30",X"50",X"D4",X"50",X"0C",X"F8",X"9B",X"5C",
		X"07",X"00",X"A0",X"3B",X"E8",X"60",X"18",X"70",X"38",X"50",X"D0",X"48",X"04",X"FA",X"A0",X"56",
		X"05",X"01",X"80",X"3C",X"F8",X"10",X"18",X"50",X"38",X"50",X"EC",X"50",X"C8",X"42",X"AB",X"4C",
		X"05",X"01",X"00",X"38",X"E8",X"60",X"18",X"60",X"40",X"60",X"C8",X"58",X"E8",X"04",X"AA",X"55",
		X"06",X"01",X"C0",X"37",X"E8",X"50",X"18",X"60",X"40",X"60",X"D0",X"50",X"EC",X"02",X"A9",X"5A",
		X"06",X"04",X"00",X"37",X"E8",X"50",X"18",X"60",X"40",X"60",X"F4",X"08",X"D4",X"56",X"A7",X"5C",
		X"07",X"05",X"00",X"37",X"E8",X"40",X"20",X"70",X"40",X"60",X"D8",X"58",X"F4",X"00",X"A8",X"59",
		X"05",X"03",X"80",X"39",X"E8",X"50",X"18",X"60",X"40",X"60",X"DC",X"50",X"F0",X"FE",X"AD",X"48",
		X"05",X"02",X"00",X"3B",X"F0",X"40",X"10",X"50",X"40",X"60",X"DC",X"58",X"EC",X"02",X"B1",X"3F",
		X"03",X"02",X"80",X"3E",X"00",X"10",X"18",X"50",X"38",X"60",X"FC",X"40",X"DC",X"56",X"A8",X"45",
		X"08",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"58",X"1C",X"32",X"EA",X"1F",
		X"06",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"2C",X"32",X"E7",X"20",
		X"08",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"48",X"EC",X"00",X"12",X"17",
		X"04",X"02",X"00",X"60",X"00",X"60",X"20",X"60",X"38",X"50",X"E0",X"68",X"F8",X"04",X"95",X"74",
		X"04",X"03",X"80",X"79",X"00",X"50",X"18",X"60",X"38",X"50",X"FC",X"08",X"E4",X"60",X"9F",X"69",
		X"03",X"03",X"00",X"81",X"00",X"40",X"18",X"60",X"30",X"40",X"F8",X"10",X"E8",X"5C",X"9F",X"67",
		X"04",X"02",X"80",X"85",X"00",X"50",X"20",X"60",X"38",X"50",X"EC",X"60",X"F4",X"08",X"9A",X"6E",
		X"03",X"01",X"40",X"81",X"00",X"40",X"20",X"60",X"38",X"60",X"F0",X"60",X"F4",X"04",X"A2",X"58",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"38",X"E4",X"08",X"FB",X"44",
		X"07",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"E0",X"08",X"FD",X"49",
		X"05",X"08",X"00",X"30",X"08",X"50",X"20",X"40",X"40",X"60",X"EC",X"58",X"DC",X"1E",X"A7",X"5D",
		X"04",X"08",X"00",X"2C",X"08",X"50",X"20",X"40",X"40",X"50",X"F0",X"48",X"E0",X"1C",X"A8",X"5D",
		X"05",X"08",X"00",X"2B",X"00",X"50",X"28",X"50",X"40",X"60",X"EC",X"48",X"E8",X"18",X"A7",X"5E",
		X"06",X"06",X"00",X"2B",X"00",X"50",X"20",X"40",X"38",X"50",X"F0",X"18",X"E8",X"56",X"A8",X"5D",
		X"03",X"06",X"00",X"2D",X"00",X"50",X"20",X"40",X"38",X"60",X"F0",X"18",X"E4",X"4C",X"A3",X"5F",
		X"03",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"30",X"F8",X"42",X"DD",X"6C",
		X"05",X"06",X"00",X"41",X"00",X"50",X"18",X"40",X"30",X"60",X"F8",X"10",X"E8",X"62",X"9F",X"6F",
		X"05",X"04",X"00",X"75",X"00",X"50",X"20",X"50",X"30",X"40",X"FC",X"08",X"E8",X"62",X"9F",X"6F",
		X"07",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"F8",X"1C",X"DF",X"13",
		X"02",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"F4",X"28",X"E7",X"11",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"A0",X"7C",X"08",X"70",X"20",X"60",X"38",X"60",X"FC",X"18",X"EC",X"6A",X"8E",X"71",
		X"02",X"01",X"C0",X"73",X"08",X"40",X"18",X"40",X"38",X"50",X"F4",X"48",X"DC",X"58",X"97",X"6D",
		X"02",X"01",X"C0",X"72",X"10",X"30",X"18",X"20",X"28",X"30",X"F4",X"38",X"D8",X"5C",X"99",X"6D",
		X"03",X"00",X"E0",X"79",X"18",X"40",X"28",X"30",X"10",X"10",X"F4",X"50",X"CC",X"54",X"9F",X"5E",
		X"0E",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"E0",X"53",X"10",X"50",X"08",X"00",X"38",X"60",X"00",X"58",X"C0",X"76",X"91",X"74",
		X"02",X"01",X"00",X"4D",X"08",X"60",X"18",X"60",X"38",X"60",X"FC",X"00",X"C0",X"72",X"9A",X"64",
		X"03",X"03",X"80",X"45",X"08",X"10",X"20",X"50",X"30",X"60",X"04",X"60",X"C4",X"76",X"9A",X"71",
		X"04",X"03",X"80",X"3D",X"08",X"00",X"20",X"60",X"30",X"60",X"04",X"68",X"C8",X"72",X"9E",X"71",
		X"04",X"03",X"00",X"39",X"00",X"00",X"18",X"60",X"30",X"60",X"00",X"60",X"C8",X"5E",X"A0",X"65",
		X"03",X"03",X"00",X"36",X"08",X"00",X"18",X"60",X"30",X"60",X"00",X"60",X"C4",X"64",X"9F",X"64",
		X"06",X"01",X"C0",X"35",X"18",X"60",X"28",X"50",X"08",X"00",X"00",X"58",X"B8",X"72",X"9C",X"68",
		X"04",X"01",X"C0",X"39",X"00",X"60",X"20",X"60",X"30",X"60",X"00",X"00",X"B8",X"70",X"9C",X"65",
		X"05",X"03",X"80",X"47",X"00",X"60",X"20",X"60",X"30",X"60",X"00",X"08",X"C4",X"60",X"9C",X"6C",
		X"03",X"06",X"00",X"50",X"F8",X"60",X"20",X"60",X"38",X"60",X"FC",X"08",X"D8",X"64",X"9D",X"75",
		X"04",X"07",X"00",X"53",X"F8",X"60",X"20",X"60",X"38",X"60",X"F8",X"08",X"DC",X"6A",X"9E",X"74",
		X"02",X"07",X"00",X"4F",X"F8",X"60",X"20",X"60",X"38",X"60",X"FC",X"08",X"E0",X"6A",X"9F",X"71",
		X"04",X"01",X"C0",X"43",X"F8",X"60",X"28",X"50",X"38",X"60",X"E0",X"60",X"F8",X"F6",X"9E",X"69",
		X"0E",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"40",X"F8",X"18",X"E0",X"29",
		X"03",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"48",X"F8",X"36",X"E7",X"0B",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"80",X"4E",X"00",X"50",X"28",X"50",X"38",X"60",X"E4",X"60",X"F0",X"0A",X"91",X"77",
		X"03",X"04",X"00",X"51",X"F8",X"50",X"20",X"40",X"38",X"60",X"FC",X"18",X"E0",X"5E",X"8E",X"7B",
		X"04",X"02",X"80",X"54",X"F8",X"50",X"20",X"50",X"38",X"70",X"F8",X"08",X"D0",X"5E",X"91",X"79",
		X"03",X"01",X"C0",X"51",X"00",X"60",X"28",X"60",X"40",X"70",X"C0",X"68",X"F4",X"00",X"95",X"73",
		X"03",X"01",X"40",X"4F",X"00",X"70",X"28",X"50",X"38",X"60",X"B8",X"78",X"F0",X"02",X"9A",X"6D",
		X"03",X"01",X"80",X"34",X"00",X"60",X"30",X"70",X"38",X"60",X"F4",X"08",X"BC",X"72",X"9B",X"6E",
		X"03",X"02",X"80",X"2C",X"00",X"60",X"30",X"70",X"40",X"70",X"F0",X"10",X"C4",X"6E",X"96",X"7A",
		X"04",X"05",X"00",X"2F",X"00",X"60",X"28",X"60",X"40",X"70",X"F8",X"08",X"C8",X"64",X"9A",X"71",
		X"04",X"07",X"00",X"32",X"00",X"60",X"28",X"50",X"38",X"60",X"F4",X"10",X"D4",X"64",X"A1",X"60",
		X"03",X"03",X"80",X"3E",X"F8",X"60",X"20",X"30",X"30",X"50",X"F8",X"08",X"E0",X"5C",X"A3",X"5C",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"18",X"D8",X"0E",X"E9",X"39",
		X"04",X"06",X"00",X"4F",X"F8",X"70",X"28",X"50",X"40",X"60",X"E4",X"60",X"F0",X"14",X"98",X"75",
		X"03",X"06",X"00",X"66",X"F8",X"60",X"28",X"60",X"38",X"50",X"FC",X"08",X"E8",X"5E",X"9C",X"6B",
		X"03",X"03",X"80",X"6F",X"F8",X"60",X"28",X"50",X"30",X"50",X"FC",X"00",X"EC",X"5C",X"99",X"69",
		X"17",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"80",X"74",X"08",X"40",X"18",X"50",X"30",X"50",X"FC",X"18",X"F0",X"64",X"8F",X"7A",
		X"03",X"05",X"00",X"74",X"00",X"50",X"18",X"60",X"30",X"50",X"00",X"10",X"EC",X"60",X"97",X"75",
		X"04",X"06",X"00",X"6E",X"00",X"50",X"18",X"60",X"28",X"40",X"FC",X"08",X"E8",X"60",X"A1",X"6A",
		X"04",X"05",X"00",X"74",X"00",X"50",X"18",X"60",X"28",X"40",X"F4",X"08",X"E8",X"5C",X"A3",X"68",
		X"03",X"06",X"00",X"75",X"00",X"50",X"18",X"60",X"28",X"40",X"F8",X"10",X"E4",X"5C",X"A3",X"6A",
		X"03",X"06",X"00",X"7B",X"00",X"50",X"18",X"50",X"30",X"40",X"FC",X"10",X"E4",X"60",X"A5",X"66",
		X"03",X"04",X"00",X"89",X"00",X"00",X"18",X"40",X"28",X"40",X"FC",X"58",X"E0",X"66",X"A6",X"67",
		X"03",X"00",X"C0",X"A2",X"F8",X"60",X"28",X"60",X"28",X"20",X"D8",X"60",X"F4",X"06",X"AA",X"53",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"00",X"5D",X"00",X"50",X"18",X"60",X"38",X"60",X"F8",X"20",X"EC",X"4A",X"95",X"72",
		X"03",X"06",X"00",X"6D",X"00",X"60",X"18",X"60",X"38",X"60",X"00",X"10",X"EC",X"58",X"97",X"70",
		X"03",X"04",X"00",X"72",X"00",X"60",X"18",X"40",X"30",X"50",X"E4",X"60",X"F4",X"06",X"A1",X"5F",
		X"03",X"01",X"40",X"7D",X"00",X"50",X"28",X"50",X"38",X"50",X"E0",X"58",X"E4",X"10",X"A9",X"4C",
		X"03",X"00",X"70",X"81",X"00",X"10",X"10",X"30",X"38",X"60",X"F8",X"50",X"D8",X"52",X"A1",X"52",
		X"03",X"00",X"40",X"89",X"F8",X"40",X"10",X"30",X"38",X"50",X"D0",X"48",X"04",X"F2",X"A5",X"4E",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"50",X"E8",X"36",X"CC",X"4F",
		X"07",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"48",X"F0",X"3A",X"D3",X"4B",
		X"08",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"48",X"F0",X"32",X"D7",X"3F",
		X"08",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"48",X"F0",X"30",X"D7",X"4A",
		X"09",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"48",X"F0",X"2E",X"D0",X"44",
		X"05",X"00",X"C0",X"36",X"E8",X"30",X"18",X"30",X"30",X"40",X"C8",X"58",X"F8",X"00",X"AC",X"49",
		X"05",X"00",X"C0",X"35",X"E8",X"40",X"18",X"40",X"30",X"40",X"CC",X"50",X"EC",X"FE",X"A7",X"59",
		X"04",X"01",X"40",X"30",X"F0",X"40",X"18",X"30",X"38",X"60",X"D8",X"70",X"E0",X"08",X"A5",X"6B",
		X"06",X"03",X"80",X"2E",X"F8",X"40",X"20",X"40",X"40",X"60",X"DC",X"60",X"E0",X"0C",X"AB",X"5E",
		X"08",X"07",X"00",X"30",X"00",X"60",X"10",X"10",X"40",X"70",X"E4",X"50",X"E4",X"10",X"B5",X"53",
		X"04",X"03",X"00",X"42",X"00",X"30",X"10",X"30",X"40",X"60",X"E0",X"48",X"E0",X"0C",X"B9",X"41",
		X"02",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"07",X"00",X"4E",X"00",X"60",X"28",X"30",X"38",X"60",X"F0",X"28",X"DC",X"4E",X"A5",X"60",
		X"02",X"05",X"00",X"70",X"00",X"40",X"10",X"20",X"38",X"40",X"F4",X"08",X"DC",X"58",X"AC",X"55",
		X"03",X"03",X"00",X"7E",X"F8",X"50",X"18",X"50",X"40",X"50",X"F8",X"08",X"CC",X"48",X"AC",X"50",
		X"0B",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"C0",X"7D",X"00",X"60",X"18",X"70",X"48",X"70",X"FC",X"08",X"C0",X"66",X"9F",X"69",
		X"03",X"02",X"00",X"91",X"00",X"60",X"18",X"70",X"48",X"70",X"FC",X"08",X"BC",X"66",X"A3",X"64",
		X"03",X"01",X"80",X"9C",X"00",X"60",X"18",X"60",X"40",X"60",X"F8",X"00",X"BC",X"60",X"A5",X"64",
		X"02",X"01",X"00",X"A5",X"00",X"70",X"18",X"60",X"40",X"60",X"BC",X"60",X"F8",X"00",X"A7",X"5E",
		X"03",X"01",X"00",X"B1",X"08",X"70",X"20",X"70",X"40",X"60",X"BC",X"70",X"F4",X"02",X"A6",X"5E",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"05",X"00",X"36",X"08",X"40",X"28",X"60",X"38",X"50",X"F4",X"58",X"F0",X"14",X"8E",X"7E",
		X"03",X"07",X"00",X"3A",X"08",X"50",X"28",X"60",X"38",X"50",X"F4",X"60",X"EC",X"10",X"93",X"73",
		X"05",X"06",X"00",X"39",X"00",X"50",X"28",X"50",X"38",X"50",X"F0",X"60",X"EC",X"0C",X"9C",X"67",
		X"03",X"07",X"00",X"3B",X"08",X"50",X"28",X"40",X"38",X"60",X"EC",X"60",X"E8",X"12",X"9F",X"72",
		X"03",X"06",X"00",X"3A",X"08",X"50",X"28",X"40",X"40",X"60",X"EC",X"58",X"E4",X"1C",X"A0",X"71",
		X"03",X"02",X"80",X"71",X"00",X"40",X"28",X"30",X"38",X"40",X"E8",X"68",X"E8",X"14",X"A1",X"70",
		X"1A",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"50",X"08",X"40",X"CF",X"35",
		X"03",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"58",X"1C",X"2E",X"E5",X"47",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"38",X"0C",X"42",X"E3",X"12",
		X"02",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"04",X"34",X"CD",X"24",
		X"03",X"05",X"00",X"47",X"10",X"50",X"20",X"50",X"30",X"60",X"F4",X"70",X"E8",X"1C",X"98",X"6E",
		X"04",X"06",X"00",X"3D",X"08",X"50",X"20",X"40",X"38",X"60",X"F0",X"60",X"E8",X"1A",X"9E",X"6D",
		X"05",X"06",X"00",X"32",X"00",X"50",X"20",X"40",X"38",X"50",X"F0",X"58",X"E4",X"1C",X"A4",X"6A",
		X"05",X"06",X"00",X"33",X"00",X"50",X"20",X"30",X"38",X"40",X"EC",X"50",X"E4",X"14",X"AA",X"61",
		X"03",X"06",X"00",X"39",X"00",X"50",X"18",X"20",X"40",X"50",X"E8",X"50",X"F0",X"0E",X"AB",X"66",
		X"03",X"01",X"40",X"47",X"00",X"40",X"18",X"20",X"40",X"50",X"E8",X"50",X"AC",X"60",X"DE",X"12",
		X"1A",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"60",X"00",X"34",X"D0",X"24",
		X"03",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"F0",X"FA",X"FC",X"43",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"05",X"00",X"49",X"08",X"40",X"10",X"30",X"30",X"50",X"F4",X"50",X"E4",X"16",X"9A",X"75",
		X"05",X"06",X"00",X"3D",X"00",X"30",X"10",X"50",X"40",X"50",X"F0",X"50",X"E8",X"0A",X"A1",X"6B",
		X"05",X"04",X"00",X"35",X"10",X"40",X"18",X"20",X"40",X"60",X"E8",X"58",X"A8",X"5E",X"D7",X"19",
		X"05",X"01",X"C0",X"30",X"00",X"20",X"18",X"60",X"40",X"50",X"E4",X"50",X"DC",X"0E",X"AB",X"55",
		X"03",X"01",X"40",X"35",X"F8",X"40",X"20",X"60",X"48",X"70",X"DC",X"50",X"E8",X"00",X"AA",X"46",
		X"0A",X"00",X"E0",X"2F",X"F8",X"40",X"18",X"60",X"48",X"60",X"E0",X"40",X"F4",X"02",X"93",X"65",
		X"08",X"00",X"A0",X"32",X"F0",X"40",X"18",X"60",X"30",X"40",X"DC",X"50",X"04",X"FC",X"8D",X"6E",
		X"06",X"00",X"50",X"34",X"F8",X"30",X"20",X"30",X"38",X"40",X"E4",X"38",X"F8",X"02",X"8B",X"71",
		X"06",X"00",X"70",X"35",X"08",X"10",X"20",X"40",X"38",X"50",X"F4",X"50",X"E8",X"1A",X"90",X"67",
		X"0B",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"00",X"42",X"DD",X"1F",
		X"06",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"40",X"E4",X"00",X"E7",X"42",
		X"05",X"03",X"00",X"8E",X"18",X"60",X"30",X"50",X"10",X"00",X"F0",X"58",X"E0",X"64",X"99",X"70",
		X"03",X"02",X"80",X"8A",X"18",X"60",X"08",X"00",X"28",X"50",X"EC",X"60",X"DC",X"66",X"9C",X"6B",
		X"04",X"02",X"80",X"B1",X"00",X"10",X"18",X"50",X"30",X"30",X"F0",X"58",X"DC",X"64",X"A2",X"6D",
		X"02",X"02",X"80",X"C7",X"00",X"00",X"18",X"60",X"28",X"30",X"F0",X"50",X"E0",X"5C",X"A2",X"6E",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"02",X"00",X"2D",X"08",X"70",X"20",X"50",X"40",X"50",X"C0",X"58",X"F0",X"04",X"AD",X"5B",
		X"07",X"03",X"00",X"2C",X"08",X"60",X"20",X"60",X"40",X"50",X"F8",X"08",X"BC",X"78",X"A8",X"5C",
		X"05",X"02",X"80",X"2A",X"08",X"70",X"20",X"60",X"38",X"60",X"BC",X"78",X"A4",X"66",X"F6",X"01",
		X"05",X"01",X"C0",X"27",X"00",X"60",X"20",X"60",X"38",X"60",X"C0",X"60",X"F4",X"00",X"A0",X"74",
		X"06",X"01",X"80",X"26",X"08",X"70",X"18",X"60",X"38",X"60",X"BC",X"60",X"F0",X"00",X"A0",X"76",
		X"08",X"01",X"80",X"26",X"00",X"60",X"18",X"50",X"30",X"40",X"BC",X"60",X"F4",X"00",X"9F",X"78",
		X"08",X"02",X"00",X"29",X"00",X"60",X"18",X"60",X"30",X"30",X"BC",X"70",X"04",X"FC",X"9B",X"77",
		X"06",X"01",X"80",X"2D",X"00",X"50",X"18",X"50",X"28",X"20",X"B4",X"78",X"0C",X"FC",X"9B",X"71",
		X"03",X"01",X"00",X"39",X"00",X"50",X"18",X"50",X"30",X"50",X"B4",X"60",X"F8",X"FC",X"9C",X"6D",
		X"03",X"00",X"E0",X"3E",X"00",X"40",X"18",X"50",X"30",X"50",X"B0",X"68",X"F8",X"00",X"99",X"73",
		X"03",X"01",X"40",X"50",X"00",X"60",X"18",X"50",X"28",X"50",X"B0",X"70",X"00",X"FE",X"99",X"6E",
		X"04",X"01",X"40",X"68",X"00",X"60",X"18",X"50",X"28",X"60",X"B0",X"70",X"0C",X"00",X"9A",X"69",
		X"03",X"00",X"C0",X"6D",X"00",X"60",X"18",X"60",X"20",X"40",X"B4",X"60",X"04",X"FC",X"9E",X"64",
		X"03",X"00",X"A0",X"70",X"08",X"60",X"20",X"50",X"30",X"40",X"B0",X"60",X"08",X"00",X"9C",X"65",
		X"03",X"00",X"40",X"7D",X"08",X"50",X"28",X"30",X"18",X"10",X"AC",X"70",X"10",X"02",X"9C",X"61",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"02",X"80",X"54",X"10",X"20",X"18",X"50",X"30",X"60",X"00",X"70",X"BC",X"76",X"A3",X"6C",
		X"04",X"02",X"80",X"51",X"08",X"10",X"18",X"60",X"30",X"60",X"04",X"68",X"BC",X"62",X"A0",X"72",
		X"03",X"03",X"00",X"4B",X"00",X"00",X"20",X"60",X"30",X"60",X"04",X"68",X"B8",X"6C",X"A0",X"71",
		X"05",X"02",X"80",X"43",X"00",X"70",X"20",X"60",X"28",X"40",X"B4",X"68",X"08",X"FC",X"A2",X"61",
		X"04",X"02",X"00",X"41",X"00",X"00",X"20",X"70",X"40",X"50",X"04",X"60",X"B4",X"62",X"9E",X"6C",
		X"04",X"01",X"C0",X"3F",X"00",X"60",X"20",X"60",X"40",X"50",X"FC",X"00",X"B4",X"6C",X"9B",X"71",
		X"04",X"02",X"00",X"3C",X"00",X"00",X"18",X"60",X"38",X"40",X"00",X"60",X"B4",X"6C",X"9B",X"6F",
		X"05",X"01",X"80",X"3E",X"18",X"50",X"00",X"00",X"28",X"40",X"00",X"50",X"B0",X"72",X"97",X"74",
		X"05",X"01",X"C0",X"41",X"00",X"00",X"18",X"70",X"30",X"60",X"00",X"58",X"B0",X"70",X"98",X"72",
		X"03",X"02",X"00",X"4A",X"18",X"70",X"30",X"50",X"08",X"00",X"00",X"50",X"B0",X"74",X"9B",X"67",
		X"03",X"01",X"C0",X"5A",X"18",X"60",X"10",X"00",X"28",X"50",X"FC",X"58",X"B0",X"6A",X"97",X"70",
		X"03",X"00",X"E0",X"63",X"00",X"00",X"18",X"60",X"38",X"60",X"00",X"48",X"AC",X"74",X"9E",X"62",
		X"03",X"00",X"A0",X"69",X"08",X"40",X"18",X"50",X"38",X"50",X"B4",X"68",X"F4",X"00",X"A3",X"5B",
		X"04",X"00",X"70",X"74",X"00",X"50",X"20",X"50",X"40",X"60",X"FC",X"00",X"B0",X"78",X"9D",X"64",
		X"03",X"00",X"80",X"83",X"00",X"60",X"20",X"50",X"40",X"70",X"B4",X"70",X"04",X"FE",X"9C",X"6A",
		X"02",X"00",X"38",X"88",X"00",X"50",X"20",X"60",X"40",X"60",X"B0",X"70",X"04",X"FE",X"A5",X"4B",
		X"04",X"00",X"38",X"80",X"08",X"40",X"20",X"40",X"38",X"50",X"B4",X"78",X"FC",X"FA",X"B5",X"39",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"58",X"20",X"36",X"E5",X"20",
		X"05",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"50",X"1C",X"36",X"ED",X"20",
		X"08",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"60",X"18",X"26",X"F4",X"20",
		X"06",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"50",X"1C",X"26",X"ED",X"2A",
		X"03",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"18",X"42",X"E0",X"3E",
		X"0A",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"50",X"FC",X"10",X"D0",X"5E",
		X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"03",X"00",X"34",X"F8",X"50",X"20",X"70",X"30",X"60",X"F8",X"08",X"C4",X"5A",X"95",X"78",
		X"06",X"04",X"00",X"2D",X"F8",X"50",X"20",X"60",X"28",X"40",X"F8",X"18",X"BC",X"70",X"9F",X"6D",
		X"03",X"02",X"80",X"29",X"00",X"60",X"20",X"50",X"30",X"40",X"F4",X"08",X"C0",X"64",X"9C",X"7A",
		X"05",X"01",X"40",X"26",X"00",X"60",X"20",X"70",X"38",X"50",X"C8",X"48",X"EC",X"00",X"9F",X"79",
		X"06",X"00",X"A0",X"24",X"00",X"40",X"20",X"70",X"38",X"50",X"C0",X"48",X"EC",X"02",X"A5",X"6B",
		X"09",X"00",X"70",X"20",X"00",X"40",X"20",X"70",X"38",X"40",X"C4",X"40",X"E8",X"FE",X"A5",X"6F",
		X"06",X"00",X"A0",X"23",X"00",X"40",X"20",X"60",X"38",X"40",X"B0",X"78",X"F8",X"FE",X"9F",X"79",
		X"04",X"00",X"E0",X"29",X"00",X"60",X"20",X"60",X"38",X"60",X"B4",X"68",X"F4",X"02",X"A4",X"61",
		X"06",X"01",X"40",X"32",X"00",X"60",X"20",X"60",X"40",X"60",X"FC",X"00",X"B4",X"68",X"A5",X"5F",
		X"05",X"01",X"40",X"3E",X"F8",X"60",X"20",X"60",X"38",X"60",X"B8",X"68",X"F4",X"02",X"A4",X"68",
		X"04",X"02",X"80",X"58",X"08",X"00",X"20",X"60",X"38",X"60",X"F0",X"58",X"C0",X"66",X"A5",X"69",
		X"03",X"01",X"00",X"65",X"E8",X"60",X"20",X"60",X"30",X"50",X"C4",X"60",X"FC",X"00",X"A7",X"69",
		X"03",X"01",X"40",X"6E",X"E8",X"60",X"20",X"60",X"28",X"40",X"CC",X"58",X"04",X"FC",X"A9",X"62",
		X"03",X"01",X"00",X"77",X"E8",X"50",X"20",X"60",X"28",X"30",X"D4",X"58",X"04",X"FE",X"A8",X"65",
		X"05",X"00",X"C0",X"76",X"E8",X"50",X"20",X"60",X"28",X"20",X"D8",X"58",X"00",X"FC",X"A7",X"69",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"80",X"45",X"00",X"60",X"20",X"40",X"30",X"50",X"00",X"18",X"BC",X"60",X"A1",X"65",
		X"03",X"06",X"00",X"4B",X"08",X"60",X"28",X"60",X"38",X"60",X"00",X"00",X"CC",X"6E",X"9D",X"6A",
		X"05",X"06",X"00",X"3E",X"08",X"60",X"28",X"50",X"38",X"50",X"EC",X"10",X"D4",X"5C",X"AF",X"63",
		X"05",X"06",X"00",X"38",X"00",X"50",X"20",X"30",X"38",X"40",X"EC",X"10",X"DC",X"50",X"B6",X"5D",
		X"06",X"06",X"00",X"37",X"00",X"50",X"20",X"30",X"38",X"40",X"E0",X"50",X"E4",X"16",X"BC",X"58",
		X"03",X"06",X"00",X"3E",X"00",X"50",X"20",X"30",X"38",X"50",X"E4",X"50",X"E4",X"16",X"B9",X"5B",
		X"04",X"04",X"00",X"4A",X"00",X"40",X"20",X"30",X"38",X"40",X"E4",X"48",X"B8",X"60",X"DF",X"11",
		X"05",X"02",X"00",X"6D",X"00",X"50",X"28",X"40",X"38",X"40",X"E4",X"60",X"E0",X"0C",X"BB",X"5A",
		X"05",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"38",X"F0",X"42",X"C6",X"40",
		X"05",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"40",X"F0",X"3E",X"C0",X"41",
		X"07",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"30",X"20",X"3A",X"EA",X"28",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"F8",X"34",X"D1",X"27",
		X"02",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"58",X"F0",X"FA",X"F5",X"24",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"80",X"5E",X"10",X"60",X"20",X"60",X"38",X"50",X"F0",X"60",X"F8",X"04",X"8F",X"74",
		X"03",X"01",X"80",X"4A",X"08",X"40",X"20",X"60",X"38",X"60",X"04",X"18",X"F0",X"60",X"8C",X"77",
		X"04",X"03",X"00",X"3C",X"00",X"50",X"20",X"60",X"40",X"60",X"00",X"08",X"F0",X"60",X"93",X"6B",
		X"03",X"03",X"80",X"36",X"00",X"10",X"28",X"60",X"40",X"60",X"FC",X"50",X"E8",X"58",X"97",X"65",
		X"05",X"01",X"80",X"30",X"00",X"50",X"28",X"60",X"38",X"60",X"F8",X"10",X"D8",X"52",X"9D",X"5C",
		X"06",X"00",X"C0",X"2A",X"00",X"50",X"28",X"70",X"38",X"60",X"CC",X"58",X"EC",X"08",X"A7",X"4B",
		X"06",X"00",X"70",X"2B",X"00",X"60",X"28",X"50",X"38",X"60",X"BC",X"78",X"F0",X"06",X"A3",X"52",
		X"06",X"00",X"38",X"27",X"08",X"60",X"30",X"60",X"30",X"30",X"C0",X"48",X"EC",X"02",X"A2",X"55",
		X"06",X"00",X"50",X"29",X"08",X"60",X"30",X"70",X"38",X"50",X"EC",X"08",X"B8",X"52",X"AF",X"42",
		X"04",X"00",X"60",X"2A",X"08",X"70",X"30",X"60",X"28",X"30",X"CC",X"78",X"E8",X"0A",X"9A",X"72",
		X"04",X"01",X"00",X"45",X"08",X"70",X"28",X"50",X"30",X"30",X"E0",X"68",X"EC",X"0A",X"A2",X"69",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"01",X"C0",X"51",X"10",X"60",X"20",X"30",X"40",X"60",X"EC",X"50",X"A8",X"6C",X"DF",X"13",
		X"04",X"05",X"00",X"3B",X"08",X"50",X"10",X"20",X"40",X"60",X"EC",X"48",X"E4",X"12",X"AD",X"67",
		X"07",X"05",X"00",X"33",X"08",X"50",X"18",X"30",X"40",X"50",X"E8",X"50",X"B4",X"60",X"E0",X"14",
		X"06",X"02",X"80",X"2D",X"08",X"40",X"18",X"20",X"38",X"60",X"E0",X"50",X"DC",X"1E",X"AE",X"5D",
		X"07",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"EC",X"22",X"DB",X"19",
		X"19",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"01",X"80",X"43",X"08",X"60",X"20",X"70",X"40",X"40",X"C4",X"60",X"F0",X"04",X"A4",X"77",
		X"03",X"03",X"80",X"3A",X"08",X"70",X"20",X"60",X"48",X"50",X"C0",X"60",X"F4",X"00",X"A8",X"61",
		X"04",X"02",X"00",X"35",X"08",X"60",X"20",X"70",X"48",X"50",X"F4",X"00",X"BC",X"74",X"A4",X"6F",
		X"04",X"01",X"C0",X"30",X"08",X"60",X"20",X"70",X"50",X"50",X"C4",X"60",X"E8",X"04",X"A6",X"6F",
		X"07",X"00",X"E0",X"2C",X"08",X"40",X"18",X"50",X"38",X"30",X"C0",X"60",X"E4",X"06",X"AB",X"61",
		X"06",X"01",X"00",X"2A",X"10",X"70",X"20",X"70",X"40",X"40",X"BC",X"60",X"E4",X"02",X"AA",X"5E",
		X"07",X"01",X"00",X"2E",X"08",X"60",X"20",X"70",X"38",X"50",X"C0",X"50",X"E4",X"04",X"A6",X"66",
		X"03",X"01",X"40",X"3C",X"08",X"60",X"20",X"70",X"38",X"50",X"B8",X"68",X"F0",X"00",X"A1",X"66",
		X"05",X"00",X"A0",X"55",X"08",X"60",X"20",X"60",X"40",X"50",X"B4",X"70",X"EC",X"02",X"9F",X"63",
		X"03",X"00",X"70",X"76",X"08",X"60",X"20",X"60",X"38",X"50",X"B0",X"68",X"F8",X"00",X"9C",X"66",
		X"04",X"00",X"40",X"87",X"20",X"60",X"30",X"30",X"08",X"00",X"08",X"50",X"AC",X"76",X"93",X"75",
		X"02",X"00",X"38",X"99",X"08",X"50",X"20",X"50",X"30",X"20",X"FC",X"00",X"B4",X"64",X"9B",X"6A",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"40",X"8C",X"00",X"60",X"30",X"50",X"30",X"20",X"F8",X"40",X"B8",X"36",X"CF",X"32",
		X"02",X"00",X"60",X"8A",X"00",X"60",X"28",X"50",X"40",X"60",X"F0",X"28",X"CC",X"1C",X"C0",X"49",
		X"03",X"00",X"38",X"80",X"00",X"40",X"28",X"50",X"40",X"70",X"F8",X"18",X"C4",X"22",X"B9",X"5E",
		X"02",X"01",X"C0",X"70",X"10",X"70",X"18",X"30",X"28",X"70",X"F8",X"00",X"BC",X"7A",X"AB",X"62",
		X"03",X"03",X"80",X"57",X"10",X"60",X"20",X"50",X"40",X"60",X"C4",X"68",X"B0",X"5C",X"F0",X"04",
		X"02",X"06",X"00",X"45",X"10",X"50",X"20",X"50",X"40",X"40",X"F4",X"18",X"C4",X"62",X"B5",X"55",
		X"05",X"07",X"00",X"35",X"10",X"60",X"20",X"40",X"38",X"40",X"E4",X"20",X"D0",X"52",X"BE",X"44",
		X"05",X"06",X"00",X"2F",X"10",X"50",X"18",X"30",X"38",X"50",X"DC",X"58",X"E0",X"18",X"BB",X"52",
		X"08",X"04",X"00",X"2E",X"18",X"50",X"10",X"20",X"38",X"50",X"DC",X"60",X"E0",X"12",X"BB",X"46",
		X"01",X"01",X"40",X"2F",X"00",X"10",X"18",X"60",X"40",X"50",X"DC",X"50",X"B0",X"4A",X"EB",X"07",
		X"0B",X"00",X"80",X"2E",X"F0",X"30",X"18",X"60",X"30",X"50",X"DC",X"40",X"F8",X"F0",X"AD",X"44",
		X"03",X"00",X"C0",X"31",X"F8",X"30",X"18",X"50",X"38",X"60",X"D8",X"48",X"04",X"FE",X"A3",X"51",
		X"0A",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"70",X"00",X"1A",X"E3",X"0E",
		X"04",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"58",X"18",X"36",X"E6",X"1C",
		X"09",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"48",X"1C",X"3E",X"E4",X"20",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"10",X"56",X"D9",X"26",
		X"02",X"05",X"00",X"48",X"08",X"50",X"20",X"40",X"30",X"40",X"EC",X"38",X"D8",X"5E",X"97",X"75",
		X"06",X"05",X"00",X"5E",X"18",X"50",X"28",X"50",X"20",X"20",X"E4",X"50",X"D4",X"66",X"9B",X"73",
		X"02",X"04",X"00",X"74",X"18",X"40",X"20",X"30",X"28",X"40",X"E4",X"50",X"D8",X"58",X"A0",X"6E",
		X"04",X"02",X"80",X"8B",X"18",X"40",X"18",X"20",X"38",X"50",X"E4",X"58",X"D8",X"64",X"A0",X"6D",
		X"02",X"01",X"40",X"97",X"08",X"10",X"20",X"50",X"40",X"60",X"E4",X"60",X"D4",X"5E",X"A0",X"70",
		X"03",X"01",X"40",X"A2",X"08",X"10",X"20",X"50",X"40",X"60",X"E8",X"60",X"D4",X"66",X"A0",X"74",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
